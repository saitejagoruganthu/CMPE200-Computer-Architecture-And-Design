module imem (
        input  wire [5:0]  a,
        output wire [31:0] y
    );

    reg [31:0] rom [0:63];

    initial begin
        $readmemh ("H:\\Masters\\Semester1\\CMPE200\\Assignment7\\memfile_withnops_updated2.dat", rom);
    end

    assign y = rom[a];
    
endmodule